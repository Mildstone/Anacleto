
module prova(
    input ca,
    output cca
    );
endmodule
